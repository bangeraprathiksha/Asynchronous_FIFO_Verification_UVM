`define DSIZE 8
`define no_of_trans 1


`define ASIZE 4
